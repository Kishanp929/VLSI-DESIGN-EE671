
	 --column 0--
	 arg1(0)<=r1(0);
	 arg2(0)<=r2(0);
	 
	 --column 1--
	 ha1:ha port map(r1(1),r2(1),arg1(1),arg2(2));
	 arg1(1)<=r3(1);
	 
	 --column 2--
	 ha2:ha port map(r1(2),r2(2),sum(0),carry(0));
	 fa1:fa port map(sum(0),r3(2),r4(2),arg1(2),arg2(3));
	 
	 --column 3--
	 fa2:fa port map(carry(0),r1(3),r2(3),sum(1),carry(1));
	 fa3:fa port map(sum(1),r3(3),r4(3),sum(2),carry(2));
	 ha3:ha port map(sum(2),r5(3),arg1(3),arg2(4));
	 
	 --column 4--
	 fa4:fa port map(r1(4),r2(4),carry(1),sum(3),carry(3));
	 fa5:fa port map(r3(4),r4(4),carry(2),sum(4),carry(4));
	 fa6: fa port map(r5(4),r6(4),sum(3),sum(5),carry(5));
	 ha4:ha port map(sum(4),sum(5),arg1(4),arg2(5));
	 
	 --column 5--
	 fa7:fa port map(r1(5),r2(5),carry(3),sum(6),carry(6));
	 fa8:fa port map(r3(5),r4(5),carry(4),sum(7),carry(7));
	 fa9:fa port map(r5(5),r6(5),carry(5),sum(8),carry(8));
	 fa10:fa port map(r7(5),sum(6),sum(7),sum(9),carry(9));
	 ha5:ha port map(sum(8),sum(9),arg1(5),arg2(6));
	 
	 --column 6--
	 fa11:fa port map(r1(6),r2(6),carry(6),sum(10),carry(10));
	 fa12:fa port map(r3(6),r4(6),carry(7),sum(11),carry(11));
	 fa13:fa port map(r5(6),r6(6),carry(8),sum(12),carry(12));
	 fa14:fa port map(r7(6),r8(6),carry(9),sum(13),carry(13));
	 fa15:fa port map(sum(10),sum(11),sum(12),sum(14),carry(14));
	 ha6:ha port map(sum(13),sum(14),arg1(6),arg2(7));
	 
	 --column 7--
	 fa16:fa port map(r1(7),r2(7),carry(10),sum(15),carry(15));
	 fa17:fa port map(r3(7),r4(7),carry(11),sum(16),carry(16));
	 fa18:fa port map(r5(7),r6(7),carry(12),sum(17),carry(17));
	 fa19:fa port map(r7(7),r8(7),carry(13),sum(18),carry(18));
	 fa20:fa port map(r9(7),sum(15),carry(14),sum(19),carry(19));	 
	 fa21:fa port map(sum(16),sum(17),sum(18),sum(20),carry(20));
	 ha7:ha port map(sum(19),sum(20),arg1(7),arg2(8));
	 
	 
	 
	 --column 8--
	 fa22:fa port map(r1(8),r2(8),carry(15),sum(21),carry(21);
	 fa24:fa port map(r3(8),r4(8),carry(16),sum(22),carry(22));
	 fa25:fa port map(r5(8),r6(8),carry(17),sum(23),carry(23));
	 fa26:fa port map(r7(8),r8(8),carry(18),sum(24),carry(24));
	 fa27:fa port map(r9(8),r10(8),carry(19),sum(25),carry(25));
	 fa28:fa port map(sum(21),sum(22),carry(20),sum(26),carry(26));
	 fa29:fa port map(sum(23),sum(24),sum(25),sum(27),carry(27));
	 ha8:ha port map(sum(26),sum(27),arg1(8),arg2(9));
	 
	 --column 9--
	 fa30:fa port map(r1(9),r2(9),carry(21),sum(28),carry(28));
	 fa31:fa port map(r3(9),r4(9),carry(22),sum(29),carry(29));
	 fa32:fa port map(r5(9),r6(9),carry(23),sum(30),carry(30));
	 fa33:fa port map(r7(9),r8(9),carry(24),sum(31),carry(31));
	 fa34:fa port map(r9(9),r10(9),carry(25),sum(32),carry(32));
	 fa35:fa port map(r11(9),carry(26),carry(27),sum(33),carry(33));
	 fa36:fa port map(sum(28),sum(29),sum(30),sum(34),carry(34));
	 fa37:fa port map(sum(31),sum(32),sum(33),sum(35),carry(35));
	 ha9:ha port map(sum(34),sum(35),arg1(9),arg2(10));

	 --column 10--
	 fa38:fa port map(r1(10),r2(10),carry(28),sum(36),carry(36));
	 fa39:fa port map(r3(10),r4(10),carry(29),sum(37),carry(37));
	 fa40:fa port map(r5(10),r6(10),carry(30),sum(38),carry(38));
	 fa41:fa port map(r7(10),r8(10),carry(31),sum(39),carry(39));
	 fa42:fa port map(r9(10),r10(10),carry(32),sum(40),carry(40));
	 fa43:fa port map(r11(10),r12(10),carry(33),sum(41),carry(41));
	 fa44:fa port map(sum(36),carry(34),carry(35),sum(42),carry(42));
	 fa45:fa port map(sum(37),sum(38),sum(38),sum(43),carry(43));
	 fa46:fa port map(sum(40),sum(41),sum(42),sum(44),carry(44));
	 ha10: ha port map(sum(43),sum(44),arg1(10),arg2(11));
	 
	 --column 11--
	 fa47:fa port map(r1(11),r2(11),carry(36),sum(45),carry(45));
	 fa48:fa port map(r3(11),r4(11),carry(37),sum(46),carry(46));
	 fa49:fa port map(r5(11),r6(11),carry(38),sum(47),carry(47));
	 fa50:fa port map(r7(11),r8(11),carry(39),sum(48),carry(48));
	 fa51:fa port map(r9(11),r10(11),carry(40),sum(49),carry(49));
	 fa52:fa port map(r11(11),r12(11),carry(41),sum(50),carry(50));
	 fa53:fa port map(r13(11),carry(42),carry(43),sum(51),carry(51));
	 fa54:fa port map(sum(45),sum(46),carry(44),sum(52),carry(52));
	 fa55:fa port map(sum(47),sum(48),sum(49),sum(53),carry(53));
	 fa56:fa port map(sum(50),sum(51),sum(52),sum(54),carry(54));
	 ha11:ha port map(sum(53),sum(54),arg1(11),arg2(12));

	 --column12--
	 fa57:fa port map(r1(12),r2(12),carry(45),sum(55),carry(55);
	 fa58:fa port map(r3(12),r4(12),carry(46),sum(56),carry(56));
	 fa59:fa port map(r5(12),r6(12),carry(47),sum(57),carry(57));
	 fa60:fa port map(r7(12),r8(12),carry(48),sum(58),carry(58));
	 fa61:fa port map(r9(12),r10(12),carry(49),sum(59),carry(59));
	 fa62:fa port map(r11(12),r12(12),carry(50),sum(60),carry(60));
	 fa63:fa port map(r13(12),r14(12),carry(51),sum(61),carry(61));
	 fa64:fa port map(carry(52),carry(53),carry(54),sum(62),carry(62));	 
	 fa65:fa port map(sum(55),sum(56),sum(57),sum(63),carry(63));
	 fa66:fa port map(sum(58),sum(59),sum(60),sum(64),carry(64));
	 fa67:fa port map(sum(61),sum(62),sum(63),sum(65),carry(65));
	 ha12:ha port map(sum(64),sum(65),arg1(12),arg2(13));
	 
	 --column13--
	 fa68:fa port map(r1(13),r2(13),carry(55),sum(66),carry(66));
	 fa69:fa port map(r3(13),r4(13),carry(56),sum(67),carry(67));
	 fa70:fa port map(r5(13),r6(13),carry(57),sum(68),carry(68));
	 fa71:fa port map(r7(13),r8(13),carry(58),sum(69),carry(69));
	 fa72:fa port map(r9(13),r10(13),carry(59),sum(70),carry(70));
	 fa73:fa port map(r11(13),r12(13),carry(60),sum(71),carry(71));
	 fa74:fa port map(r13(13),r14(13),carry(61),sum(72),carry(72));
	 fa75:fa port map(r15(13),carry(62),carry(63),sum(73),carry(73));
	 fa76:fa port map(sum(66),sum(67),carry(64),sum(74),carry(74));
	 fa77:fa port map(sum(68),sum(69),carry(65),sum(75),carry(75));
	 fa78:fa port map(sum(70),sum(71),sum(72),sum(76),carry(76));
	 fa79:fa port map(sum(73),sum(74),sum(75),sum(77),carry(77));
	 ha13:ha port map(sum(76),sum(77),arg1(13),arg2(14));
	 
	 --column 14--
	 fa80:fa port map(r1(14),r2(14),carry(66),sum(78),carry(78));
	 fa81:fa port map(r3(14),r4(14),carry(67),sum(79),carry(79));
	 fa82:fa port map(r5(14),r6(14),carry(68),sum(80),carry(80));
	 fa83:fa port map(r7(14),r8(14),carry(69),sum(81),carry(81));
	 fa84:fa port map(r9(14),r10(14),carry(70),sum(82),carry(82));
	 fa85:fa port map(r11(14),r12(14),carry(71),sum(83),carry(83));
	 fa86:fa port map(r13(14),r14(14),carry(72),sum(84),carry(84));
	 fa87:fa port map(r15(14),r16(14),carry(73),sum(85),carry(85));
	 fa88:fa port map(carry(74),carry(75),carry(76),sum(86),carry(86));
	 fa89:fa port map(sum(78),sum(79),carry(77),sum(87),carry(87));
	 fa90:fa port map(sum(80),sum(81),sum(82),sum(88),carry(88));
	 fa91:fa port map(sum(83),sum(84),sum(85),sum(89),carry(89));
	 fa92:fa port map(sum(86),sum(87),sum(88),sum(90),carry(90));
	 ha14:ha port map(sum(89),sum(90),arg1(14),arg2(15));
	 
	 --column 15--
	 fa93:fa port map(r1(15),r2(15),carry(78),sum(91),carry(91));
	 fa94:fa port map(r3(15),r4(15),carry(79),sum(92),carry(92));
	 fa95:fa port map(r5(15),r6(15),carry(80),sum(93),carry(93));
	 fa96:fa port map(r7(15),r8(15),carry(81),sum(94),carry(94));
	 fa97:fa port map(r9(15),r10(15),carry(82),sum(95),carry(95));
	 fa98:fa port map(r11(15),r12(15),carry(83),sum(96),carry(96));
	 fa99:fa port map(r13(15),r14(15),carry(84),sum(97),carry(97));
	 fa100:fa port map(r15(15),r16(15),carry(85),sum(98),carry(98));
	 fa101:fa port map(r17(17),carry(86),carry(87),sum(99),carry(99));
	 fa102:fa port map(carry(88),carry(89),carry(90),sum(100),carry(100));
	 fa103:fa port map(sum(91),sum(92),sum(93),sum(101),carry(101));
	 fa104:fa port map(sum(94),sum(95),sum(96),sum(102),carry(102));
	 fa105:fa port map(sum(97),sum(98),sum(99),sum(103),sum(103));
	 fa106:fa port map(sum(100),sum(101),sum(102),sum(104),carry(104));
	 ha15:ha port map(sum(103),sum(104),arg1(15),arg2(16));
	 
	 --column 16--  16-15 rows after r1 are 0
	 fa107:fa port map(r1(16),r3(16),carry(91),sum(105),carry(105));
	 fa108:fa port map(r4(16),r5(16),carry(92),sum(106),carry(106));
	 fa109:fa port map(r6(16),r7(16),carry(93),sum(107),carry(107));
	 fa110:fa port map(r8(16),r9(16),carry(94),sum(108),carry(108));
	 fa111:fa port map(r10(16),r11(16),carry(95),sum(109),carry(109));
	 fa112:fa port map(r12(16),r13(16),carry(96),sum(110),carry(110));
	 fa113:fa port map(r14(16),r15(16),carry(97),sum(111),carry(111));
	 fa114:fa port map(r16(16),r17(16),carry(98),sum(112),carry(112));
	 fa115:fa port map(carry(99),carry(100),carry(101),sum(113),carry(113));
	 fa116:fa port map(carry(102),carry(103),carry(104),sum(114),carry(114));
	 fa117:fa port map(sum(105),sum(106),sum(107),sum(115),carry(115));
	 fa118:fa port map(sum(108),sum(109),sum(110),sum(116),carry(116));
	 fa119:fa port map(sum(111),sum(112),sum(113),sum(117),carry(117));
	 fa120:fa port map(sum(114),sum(115),sum(116),sum(118),carry(118));
	 ha16:ha port map(sum(117),sum(118),arg1(16),arg2(17));
	 
	 --cloumn 17-- 2 rows are zero
	 fa121: fa port map(r1(17),r4(17),carry(105),sum(119),carry(119));
	 fa122: fa port map(r5(17),r6(17),carry(106),sum(120),carry(120));
	 fa123: fa port map(r7(17),r8(17),carry(107),sum(121),carry(121));
	 fa124: fa port map(r9(17),r10(17),carry(108),sum(122),carry(122));
	 fa125: fa port map(r11(17),r12(17),carry(109),sum(123),carry(123));
	 fa126: fa port map(r13(17),r14(17),carry(110),sum(124),carry(124));
	 fa127: fa port map(r15(17),r16(17),carry(111),sum(125),carry(125));
	 fa128: fa port map(r17(17),sum(99),sum(112),sum(126),carry(126));
	 fa129:fa port map(carry(113),carry(114),carry(115),sum(127),carry(127));
	 fa130:fa port map(carry(116),carry(117),carry(118),sum(128),carry(128));
	 fa131: fa port map(sum(119),sum(120),sum(121),sum(129),carry(129));
	 fa132: fa port map(sum(122),sum(123),sum(124),sum(130),carry(130));
	 fa133: fa port map(sum(125),sum(126),sum(127),sum(131),carry(131));
	 fa134: fa port map(sum(128),sum(129),sum(130),sum(132),carry(132));	 
	 ha17:ha port map(sum(131),sum(132),arg1(17),arg2(18));
	 
	 --cloumn 18-- 3 rows are zero
	 fa135:fa port map(r1(18),r5(18),carry(119),sum(133),carry(133));
	 fa136:fa port map(r6(18),r7(18),carry(120),sum(134),carry(134));
	 fa137:fa port map(r8(18),r9(18),carry(121),sum(135),carry(135));
	 fa138:fa port map(r10(18),r11(18),carry(122),sum(136),carry(136));
	 fa139:fa port map(r12(18),r13(18),carry(123),sum(137),carry(137));
	 fa140:fa port map(r14(18),r15(18),carry(124),sum(138),carry(138));
	 fa141:fa port map(r16(18),r17(18),carry(125),sum(139),carry(139));
	 fa142:fa port map(carry(126),carry(127),carry(128),sum(140),carry(140));
	 fa143:fa port map(carry(129),carry(130),carry(131),sum(141),carry(141));
	 fa144:fa port map(sum(133),sum(134),carry(132),sum(142),carry(142));
	 fa145:fa port map(sum(135),sum(136),sum(137),sum(143),carry(143));
	 fa146:fa port map(carry(138),carry(139),carry(140),sum(144),carry(144));
	 fa147:fa port map(carry(141),carry(142),carry(143),sum(145),carry(145));
	 ha18:ha port map(sum(144),sum(145),arg1(18),arg2(19));
	 
	 --cloumn 19-- 4 rows are zero
	 fa148:fa port map(r1(19),r6(19),carry(133),sum(146),carry(146));
	 fa149:fa port map(r7(19),r8(19),carry(134),sum(147),carry(147));
	 fa150:fa port map(r9(19),r10(19),carry(135),sum(148),carry(148));
	 fa151:fa port map(r11(19),r12(19),carry(136),sum(149),carry(149));
	 fa152:fa port map(r13(19),r14(179),carry(137),sum(150),carry(150));
	 fa153:fa port map(r15(19),r16(19),carry(138),sum(151),carry(151));
	 fa154:fa port map(r17(19),carry(139),carry(140),sum(152),carry(152));
	 fa155:fa port map(carry(141),carry(142),carry(143),sum(153),carry(153));
	 fa156:fa port map(carry(144),carry(145),sum(146),sum(154),carry(154));
	 fa157:fa port map(sum(147),sum(148),sum(149),sum(155),carry(155));
	 fa158:fa port map(sum(150),sum(151),sum(152),sum(156),carry(156));
	 fa159:fa port map(sum(153),sum(154),sum(155),sum(157),carry(157));
	 ha19:ha port map(sum(156),sum(157),arg1(19),arg2(20));
	 
	 --clomun 20 -- 5 rows are zero
	 fa160:fa port map(r1(20),r7(20),carry(146),sum(158),carry(158));
	 fa161:fa port map(r8(20),r9(20),carry(147),sum(159),carry(159));
	 fa162:fa port map(r10(20),r11(20),carry(148),sum(160),carry(160));
	 fa163:fa port map(r12(20),r13(20),carry(149),sum(161),carry(161));
	 fa164:fa port map(r14(20),r15(20),carry(150),sum(162),carry(162));
	 fa165:fa port map(r16(20),r17(20),carry(151),sum(163),carry(163));
	 fa166:fa port map(carry(152),carry(153),carry(154),sum(164),carry(164));
	 fa167:fa port map(carry(155),carry(156),carry(157),sum(165),carry(165));
	 fa168:fa port map(sum(158),sum(159),sum(160),sum(166),carry(166));
	 fa169:fa port map(sum(161),sum(162),sum(163),sum(167),carry(167));
	 fa170:fa port map(sum(164),sum(165),sum(166),sum(168),carry(168));
	 ha20:ha port map(sum(167),sum(168),arg1(20),arg2(21));
	 
	 --cloumn 21 --6 rows are zero
	 fa171:fa port map(r1(21),r8(21),carry(158),sum(169),carry(169));
	 fa172:fa port map(r9(21),r10(21),carry(159),sum(170),carry(170));
	 fa173:fa port map(r11(21),r12(21),carry(160),sum(171),carry(171));
	 fa174:fa port map(r13(21),r14(21),carry(161),sum(172),carry(172));
	 fa175:fa port map(r15(21),r16(21),carry(162),sum(173),carry(173));
	 fa176:fa port map(r17(21),carry(163),carry(164),sum(174),carry(174));
	 fa177:fa port map(carry(165),carry(166),carry(167),sum(175),carry(175));	 
	 fa178:fa port map(carry(168),sum(169),sum(170),sum(176),carry(176));
	 fa179:fa port map(sum(171),sum(172),sum(173),sum(177),carry(177));
	 fa180:fa port map(sum(174),sum(175),sum(176),sum(178),carry(178));
	 ha21:ha port map(sum(177),sum(178),arg1(21),arg2(22));

	 --clolumn 22 
	 fa181:fa port map(r1(22),r9(22),carry(169),sum(179),carry(179));
	 fa182:fa port map(r10(22),r11(22),carry(170),sum(180),carry(180));
	 fa183:fa port map(r12(22),r13(22),carry(171),sum(181),carry(181));
	 fa184:fa port map(r14(22),r15(22),carry(172),sum(182),carry(182));
	 fa185:fa port map(r16(22),r17(22),carry(173),sum(183),carry(183));
	 fa186:fa port map(carry(174),carry(175),carry(176),sum(184),carry(184));	 
	 fa187:fa port map(carry(177),carry(178)sum(179),sum(185),carry(185));
	 fa188:fa port map(sum(180),sum(181),sum(182),sum(186),carry(186));
	 fa189:fa port map(sum(183),sum(184),sum(185),sum(187),carry(187));
	 ha22:ha port map(sum(186),sum(187),arg1(22),arg2(23));	 
	 
	 --cloumn 23
	 fa190:fa port map(r1(23),r10(23),carry(179),sum(188),carry(188));
	 fa191:fa port map(r11(22),r12(23),carry(180),sum(189),carry(189));
	 fa192:fa port map(r13(22),r14(23),carry(181),sum(190),carry(190));
	 fa193:fa port map(r15(22),r16(23),carry(182),sum(191),carry(191));
	 fa194:fa port map(r17(22),carry(183),carry(184),sum(192),carry(192));
	 fa195:fa port map(carry(185),carry(186),carry(187),sum(193),carry(193));
	 fa196:fa port map(sum(188),sum(189),sum(190),sum(194),carry(194));
	 fa197:fa port map(sum(191),sum(192),sum(193),sum(195),carry(195));
	 ha23:ha port map(sum(194),sum(195),arg1(23),arg2(24));	 	 
	 
	 --column 24
	 fa198:fa port map(r1(24),r11(24),carry(188),sum(196),carry(196));
	 fa199:fa port map(r12(24),r13(24),carry(189),sum(197),carry(197));
	 fa200:fa port map(r14(24),r15(24),carry(190),sum(198),carry(198));
	 fa201:fa port map(r16(24),r17(24),carry(191),sum(199),carry(199));
	 fa202:fa port map(carry(192),carry(193),carry(194),sum(200),carry(200));
	 fa203:fa port map(carry(195),sum(196),sum(197),sum(201),carry(201));
	 fa204:fa port map(sum(198),sum(199),sum(200),sum(202),carry(202));
	 ha24:ha port map(sum(201),sum(202),arg1(24),arg2(25));
	 
	 --column 25
	 fa205:fa port map(r1(25),r12(25),carry(196),sum(203),carry(203));
	 fa206:fa port map(r13(25),r14(25),carry(197),sum(204),carry(204));
	 fa207:fa port map(r15(25),r16(25),carry(198),sum(205),carry(205));
	 fa208:fa port map(r17(25),carry(199),carry(200),sum(206),carry(206));
	 fa209:fa port map(carry(201),carry(202),sum(203),sum(207),sum(207));
	 fa210:fa port map(sum(204),sum(205),sum(206),sum(208),carry(208));
	 ha25:ha port map(sum(207),sum(208),arg1(25),arg2(26));
	 
	 --column 26
	 fa211:fa port map(r1(26),r13(26),carry(203),sum(209),carry(209));
	 fa212:fa port map(r14(26),r15(26),carry(204),sum(210),carry(210));
	 fa213:fa port map(r16(26),r17(26),carry(205),sum(211),carry(211));
	 fa214:fa port map(carry(206),carry(207),carry(208),sum(212),carry(212));
	 fa215:fa port map(sum(209),sum(210),sum(211),sum(213),carry(213));
	 ha26:ha port map(sum(212),sum(213),arg1(26),arg2(27));
	 
	 --column 27
	 fa216:fa port map(r1(27),r14(27),carry(209),sum(214),carry(214));
	 fa217:fa port map(r15(27),r16(27),carry(210),sum(215),carry(215));
	 fa218:fa port map(r17(27),carry(211),carry(212),sum(216),carry(216));
	 fa219:fa port map(carry(213),sum(214),sum(215),sum(217),carry(217));
	 ha27:ha port map(sum(216),sum(217),arg1(27),arg2(28));
	 
	 --column 28
	 fa220:fa port map(r1(28),r15(28),carry(214),sum(218),carry(218));
	 fa221:fa port map(r16(28),r17(28),carry(215),sum(219),carry(219));
	 fa222:fa port map(carry(216),carry(217),sum(218),sum(220),carry(220));
	 ha28:ha port map(sum(219),sum(220),arg1(28),arg2(29));
	 
	 --column 29
	 fa223:fa port map(r1(29),r16(29),carry(218),sum(221),carry(221));
	 fa224:fa port map(r17(29),carry(219),carry(220),sum(222),carry(222));
	 ha29:ha port map(sum(221),sum(222),arg1(29),arg2(30));
	 
	 --column 30
	 fa225:fa port map(r1(30),r17(30),carry(221),sum(223),carry(223));
	 ha30:ha port map(carry(222),sum(223),arg1(30),arg2(31));
	 
	 --column 31
	 arg1(31)<=carry(223);
	 
	 
	 
	 
	 
	 
	 





